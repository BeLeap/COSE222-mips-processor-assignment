module memory(
    input [31:0] addr, write_data,
    input MemWrite, MemRead,
    output [31:0] read_data
    );

endmodule