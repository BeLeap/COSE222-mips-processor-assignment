module control(
    input wire [6:0] inst,
    output wire RegDst, Jump, Branch, MemRead, MemToReg, ALUOp, MemWrite, ALUSrc, RegWrite
    );

endmodule