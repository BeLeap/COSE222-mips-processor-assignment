module memory(
    input wire rst, clk,
    input wire [31:0] addr, write_data,
    input wire MemWrite, MemRead,
    output wire [31:0] read_data
    );

    reg [31:0] mem [0:63];

    always @(negedge rst or posedge clk) begin
        if (!rst) begin
            mem [0] <= 32'b00000000000000000000000000000000;
            mem [1] <= 32'b00000000000000000000000000000001;
            mem [2] <= 32'b00000000000000000000000000000010;
            mem [3] <= 32'b00000000000000000000000000000011;
            mem [4] <= 32'b00000000000000000000000000000100;
            mem [5] <= 32'b00000000000000000000000000000111;
            mem [6] <= 32'b00000000000000000000000000000110;
            mem [7] <= 32'b00000000000000000000000000000111;
            mem [8] <= 32'b00000000000000000000000000001000;
            mem [9] <= 32'b00000000000000000000000000001001;
            mem [10] <= 32'b00000000000000000000000000001010;
            mem [11] <= 32'b00000000000000000000000000001011;
            mem [12] <= 32'b00000000000000000000000000001100;
            mem [13] <= 32'b00000000000000000000000000001101;
            mem [14] <= 32'b00000000000000000000000000001110;
            mem [15] <= 32'b00000000000000000000000000001111;
            mem [16] <= 32'b00000000000000000000000000010000;
            mem [17] <= 32'b00000000000000000000000000010001;
            mem [18] <= 32'b00000000000000000000000000010010;
            mem [19] <= 32'b00000000000000000000000000010011;
            mem [20] <= 32'b00000000000000000000000000010100;
            mem [21] <= 32'b00000000000000000000000000010101;
            mem [22] <= 32'b00000000000000000000000000010110;
            mem [23] <= 32'b00000000000000000000000000010111;
            mem [24] <= 32'b00000000000000000000000000011000;
            mem [25] <= 32'b00000000000000000000000000011001;
            mem [26] <= 32'b00000000000000000000000000011010;
            mem [27] <= 32'b00000000000000000000000000011011;
            mem [28] <= 32'b00000000000000000000000000011100;
            mem [29] <= 32'b00000000000000000000000000011101;
            mem [30] <= 32'b00000000000000000000000000011110;
            mem [31] <= 32'b00000000000000000000000000011111;
            mem [32] <= 32'b00000000000000000000000000000000;
            mem [33] <= 32'b00000000000000000000000000000001;
            mem [34] <= 32'b00000000000000000000000000000010;
            mem [35] <= 32'b00000000000000000000000000000011;
            mem [36] <= 32'b00000000000000000000000000000100;
            mem [37] <= 32'b00000000000000000000000000000101;
            mem [38] <= 32'b00000000000000000000000000000110;
            mem [39] <= 32'b00000000000000000000000000000111;
            mem [40] <= 32'b00000000000000000000000000001000;
            mem [41] <= 32'b00000000000000000000000000001001;
            mem [42] <= 32'b00000000000000000000000000001010;
            mem [43] <= 32'b00000000000000000000000000001011;
            mem [44] <= 32'b00000000000000000000000000001100;
            mem [45] <= 32'b00000000000000000000000000001101;
            mem [46] <= 32'b00000000000000000000000000001110;
            mem [47] <= 32'b00000000000000000000000000001111;
            mem [48] <= 32'b00000000000000000000000000010000;
            mem [49] <= 32'b00000000000000000000000000010001;
            mem [50] <= 32'b00000000000000000000000000010010;
            mem [51] <= 32'b00000000000000000000000000010011;
            mem [52] <= 32'b00000000000000000000000000010100;
            mem [53] <= 32'b00000000000000000000000000010101;
            mem [54] <= 32'b00000000000000000000000000010110;
            mem [55] <= 32'b00000000000000000000000000010111;
            mem [56] <= 32'b00000000000000000000000000011000;
            mem [57] <= 32'b00000000000000000000000000011001;
            mem [58] <= 32'b00000000000000000000000000011010;
            mem [59] <= 32'b00000000000000000000000000011011;
            mem [60] <= 32'b00000000000000000000000000011100;
            mem [61] <= 32'b00000000000000000000000000011101;
            mem [62] <= 32'b00000000000000000000000000011110;
            mem [63] <= 32'b00000000000000000000000000011111;
        end
        else if (MemWrite) begin
                mem[addr] <= write_data;
        end
    end

    assign read_data = MemWrite ? write_data : mem[addr][31:0];

endmodule